`timescale 1ns/1ps

module cpu (
    input logic clk,
    input logic rst_n
);

endmodule